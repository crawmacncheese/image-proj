*SPICE Netlist for circuit 0


.OP
.END

