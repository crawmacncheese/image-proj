*SPICE Netlist for circuit 0
M1 4 5 4 4 MMOS W=1u L=1u
M3 4 6 4 4 MMOS W=1u L=1u
M2 5 1 7 7 MMOS W=1u L=1u
M4 7 8 6 6 MMOS W=1u L=1u
M6 9 10 8 8 MMOS W=1u L=1u
M5 11 9 2 2 MMOS W=1u L=1u
M7 10 11 11 MMOS W=1u L=1u

.OP
.END

